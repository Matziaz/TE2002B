-- Encryptor