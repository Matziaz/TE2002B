----------------------------------------------------------------------------------
-- Company:		ITESM - IRS 2025
-- Author:           	Dalila Fonseca, Santiago Gonzáles, Victoria Robles, Angelo Segura
-- Create Date: 	22/04/2025
-- Design Name: 	Shift Rows
-- Module Name:		Shift Rows Module
-- Target Devices: 	DE10-Lite
-- Description: 	Shift Rows AES - Module
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity ShiftRows is
  port (
    Clk    : in     std_logic;
    Enable : in     std_logic;
    Finish : out    std_logic;
    Rst    : in     std_logic;
    TxtIn  : in     std_logic_vector(127 downto 0);
    TxtOut : out    std_logic_vector(127 downto 0)
  );
end entity ShiftRows;

architecture rtl of ShiftRows is
    -- State machine
	 type state_type is (St0, St1, St2);
	 signal present_state, next_state : state_type;
    
	 -- 16-byte arrays for input and output
	 type byte_array is array (0 to 15) of std_logic_vector(7 downto 0);
    
    signal input_bytes  : byte_array;
    signal output_bytes : byte_array;
    signal result       : std_logic_vector(127 downto 0) := (others => '0');
	 signal result_reg   : std_logic_vector(127 downto 0) := (others => '0');
    signal done         : std_logic := '0';
    signal enable_reg   : std_logic := '0';
begin

    -- Clock proces: handles state transitions
    process(Clk, Rst)
    begin
        if Rst = '1' then
				present_state <= St0;
            done <= '0';
            enable_reg <= '0';
        elsif rising_edge(Clk) then
				present_state <= next_state;
            enable_reg <= Enable;
				
				case present_state is
					when St0 =>
						done <= '0';
					when St1 =>
						-- Save processed result
						result_reg <= result;
					when St2 =>
						done <= '1';
				end case;
        end if;
    end process;
	 
	 --Next stage logic
	 process(present_state, Enable)
	 begin
		next_state <= present_state;
		
		case present_state is 
			when St0 =>
				if Enable = '1' then
					next_state <= St1;
				end if;
			when St1 =>
				next_state <= St2;
			when St2 =>
				if Enable = '0' then
					next_state <= St0;
				end if;
		end case;
	end process;
					

    -- Input separation process (combinational)
	 --Split 128-bit input into 16 bytes
    process (TxtIn)
    begin
        for i in 0 to 15 loop
            input_bytes(i) <= TxtIn(127 - i*8 downto 120 - i*8);
        end loop;
    end process;

    -- ShiftRows operation process (combinational)
    process (input_bytes)
    begin
		  -- Row 0 (no shift)	
        output_bytes(0)  <= input_bytes(0);
        output_bytes(4)  <= input_bytes(4);
        output_bytes(8)  <= input_bytes(8);
        output_bytes(12) <= input_bytes(12);
		  
		  --Row 1 (shift left by 1)
        output_bytes(1)  <= input_bytes(5);
        output_bytes(5)  <= input_bytes(9);
        output_bytes(9)  <= input_bytes(13);
        output_bytes(13) <= input_bytes(1);

		  --Row 2 (shift left by 2)
        output_bytes(2)  <= input_bytes(10);
        output_bytes(6)  <= input_bytes(14);
        output_bytes(10) <= input_bytes(2);
        output_bytes(14) <= input_bytes(6);

		  --Row 3 (shift left by 3)
        output_bytes(3)  <= input_bytes(15);
        output_bytes(7)  <= input_bytes(3);
        output_bytes(11) <= input_bytes(7);
        output_bytes(15) <= input_bytes(11);
    end process;

    -- Output reconstruction process (combinational)
	 -- Combine output bytes into 128-bit vector
    process (output_bytes)
    begin
        result <=
            output_bytes(0)  & output_bytes(1)  & output_bytes(2)  & output_bytes(3)  &
            output_bytes(4)  & output_bytes(5)  & output_bytes(6)  & output_bytes(7)  &
            output_bytes(8)  & output_bytes(9)  & output_bytes(10) & output_bytes(11) &
            output_bytes(12) & output_bytes(13) & output_bytes(14) & output_bytes(15);
	 end process;

    -- Output assignments
    TxtOut <= result_reg;
    Finish <= done;
  end architecture rtl; -- of ShiftRows

