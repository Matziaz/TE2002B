-- Decryptor