----------------------------------------------------------------------------------
-- Company:		ITESM - IRS 2025
-- Author:           	Emiliano Camacho, Obiel Rangel, Evan Santana, Alfredo Soto 
-- Create Date: 	22/04/2025
-- Design Name: 	Add Round Key
-- Module Name:		Add Round Key Module
-- Target Devices: 	DE10-Lite
-- Description: 	Add Round Key AES - Module
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity AddRoundKey is
    Port ( KeyIn  : in  STD_LOGIC_VECTOR (127 downto 0);        -- Clave de ronda
           Clk    : in     std_logic;                           --Señal de reloj
			  Enable : in     std_logic;                           --Habilita el funcionamiento
		     Rst    : in     std_logic;                           --Señal de reset  
			  TxtIn  : in     std_logic_vector(127 downto 0);      --Texto de entrada de datos de 128 bits
			  TxtOut : out    std_logic_vector(127 downto 0);     -- Texto de salida de datos de 128 bits
			  Finish : out    STD_LOGIC:='0');                     --Indica fin de funcionamiento
end AddRoundKey;

architecture Behavioral of AddRoundKey is
   -- Señales intermedias para almacenar entradas
	signal cipher : STD_LOGIC_VECTOR (127 downto 0);
	signal round : STD_LOGIC_VECTOR (127 downto 0);
	
	 -- Tipo de dato para almacenamiento byte a byte
	type tipo_SRAM is ARRAY (0 to 15) of STD_LOGIC_VECTOR (7 downto 0);
	
	-- Memoria para almacenar texto y clave por bytes
	signal memoria_cipher : tipo_SRAM;
	signal memoria_key : tipo_SRAM;
	
	-- Señal de control interna para Finish
	signal Flag: STD_LOGIC := '0';
	
	
begin
	cipher <= TxtIn;
	round <= KeyIn;
	
	-- Proceso principal: AddRoundKey
	process(Clk,Enable)
	begin
	if (rising_edge(Clk) and Enable = '1')then
	-- División del texto de entrada en 16 bytes (128 bits total)
   memoria_cipher(0) <= cipher(7 downto 0);
	memoria_cipher(1) <= cipher(15 downto 8);
	memoria_cipher(2) <= cipher(23 downto 16);
	memoria_cipher(3) <= cipher(31 downto 24);
	memoria_cipher(4) <= cipher(39 downto 32);
	memoria_cipher(5) <= cipher(47 downto 40);
	memoria_cipher(6) <= cipher(55 downto 48);
	memoria_cipher(7) <= cipher(63 downto 56);
	memoria_cipher(8) <= cipher(71 downto 64);
	memoria_cipher(9) <= cipher(79 downto 72);
	memoria_cipher(10) <= cipher(87 downto 80);
	memoria_cipher(11) <= cipher(95 downto 88);
	memoria_cipher(12) <= cipher(103 downto 96);
	memoria_cipher(13) <= cipher(111 downto 104);
	memoria_cipher(14) <= cipher(119 downto 112);
	memoria_cipher(15) <= cipher(127 downto 120);
	
	-- División de la clave en 16 bytes (128 bits total)
	memoria_key(0) <= round(7 downto 0);
	memoria_key(1) <= round(15 downto 8);
	memoria_key(2) <= round(23 downto 16);
	memoria_key(3) <= round(31 downto 24);
	memoria_key(4) <= round(39 downto 32);
	memoria_key(5) <= round(47 downto 40);
	memoria_key(6) <= round(55 downto 48);
	memoria_key(7) <= round(63 downto 56);
	memoria_key(8) <= round(71 downto 64);
	memoria_key(9) <= round(79 downto 72);
	memoria_key(10) <= round(87 downto 80);
	memoria_key(11) <= round(95 downto 88);
	memoria_key(12) <= round(103 downto 96);
	memoria_key(13) <= round(111 downto 104);
	memoria_key(14) <= round(119 downto 112);
	memoria_key(15) <= round(127 downto 120);

	-- Operación XOR byte a byte
	TxtOut (7 downto 0)  <= memoria_cipher(0) xor memoria_key(0);
	TxtOut (15 downto 8) <= memoria_cipher(1) xor memoria_key(1);
	TxtOut (23 downto 16) <= memoria_cipher(2) xor memoria_key(2);
	TxtOut (31 downto 24) <= memoria_cipher(3) xor memoria_key(3);
	TxtOut (39 downto 32) <= memoria_cipher(4) xor memoria_key(4);
	TxtOut (47 downto 40) <= memoria_cipher(5) xor memoria_key(5);
	TxtOut (55 downto 48) <= memoria_cipher(6) xor memoria_key(6);
	TxtOut (63 downto 56) <= memoria_cipher(7) xor memoria_key(7);
	TxtOut (71 downto 64) <= memoria_cipher(8) xor memoria_key(8);
	TxtOut (79 downto 72) <= memoria_cipher(9) xor memoria_key(9);
	TxtOut (87 downto 80) <= memoria_cipher(10) xor memoria_key(10);
	TxtOut (95 downto 88) <= memoria_cipher(11) xor memoria_key(11);
	TxtOut (103 downto 96) <= memoria_cipher(12) xor memoria_key(12);
	TxtOut (111 downto 104) <= memoria_cipher(13) xor memoria_key(13);
	TxtOut (119 downto 112) <= memoria_cipher(14) xor memoria_key(14);
	TxtOut (127 downto 120) <= memoria_cipher(15) xor memoria_key(15);   
	end if;

	end process;	

	 -- Proceso de control: Generación de señal Finish
	process(Rst,Clk,Enable)
		 
		variable cta : STD_LOGIC_VECTOR (1 downto 0):="00";
		begin
			if Rst = '1' then
				cta := "00";
			elsif rising_edge(Clk) then
				if Enable = '1' then
				-- Incrementa contador solo si Enable está activo
					cta := cta + 1;
					-- Después de 3 ciclos (contando desde 0), activa Finish
					if cta = "11" then --2do. clock
						Flag <= '1';
					end if;
				end if;
				-- Autolimpieza de la señal Flag
				if Flag = '1' then
					Flag<='0';
				end if;
			end if;

		end process;
		
	-- Asignación de la señal interna Flag a la salida Finish
	Finish <= Flag;



end Behavioral;
